--Este Mux32_a_1 utiliza la misma logica que cualquier otro mux, con ladiferencia que tienen 32 entradas, y 32 salidas.
--Mientras que su S es de 5 bits.

library IEEE;
use IEEE.std_logic_1164.all;

entity Mux_32_a_1_21Bits is
	port (
	A, B, C, D, E, F, G, H, I, J,
	K, L, M, N, O, P, Q, R, Si, T,
	U, W, X, Y, Z, A1, B1, C1, D1, E1,
	F1, G1: in std_logic_vector (20 downto 0);
	S: in std_logic_vector (4 downto 0);
	Rout: out std_logic_vector (20 downto 0));
end Mux_32_a_1_21Bits;
 
architecture Mux_32_a_1_21Bits of Mux_32_a_1_21Bits is
component Mux32_a_1 
	port (
	a, b, c, d, e, f, g, h, i, j,
	k, l, m, n, o, p, q, r, si, t,
	u, w, x, y, z, a1, b1, c1, d1, e1,
	f1, g1: in std_logic;
	S: in std_logic_vector (4 downto 0);
	Rout: out std_logic);
end component; 

begin
	Mux_32_a_18Bits_0: Mux32_a_1 port map (A(0), B(0), C(0), D(0), E(0), F(0), G(0), H(0), I(0), J(0),
	K(0), L(0), M(0), N(0), O(0), P(0), Q(0), R(0), Si(0), T(0), U(0), W(0), X(0), Y(0), Z(0),
	A1(0), B1(0), C1(0), D1(0), E1(0), F1(0), G1(0), S, Rout(0));
	Mux_32_a_18Bits_1: Mux32_a_1 port map (A(1), B(1), C(1), D(1), E(1), F(1), G(1), H(1), I(1), J(1),
	K(1), L(1), M(1), N(1), O(1), P(1), Q(1), R(1), Si(1), T(1), U(1), W(1), X(1), Y(1), Z(1),
	A1(1), B1(1), C1(1), D1(1), E1(1), F1(1), G1(1), S, Rout(1));
	Mux_32_a_18Bits_2: Mux32_a_1 port map (A(2), B(2), C(2), D(2), E(2), F(2), G(2), H(2), I(2), J(2),
	K(2), L(2), M(2), N(2), O(2), P(2), Q(2), R(2), Si(2), T(2), U(2), W(2), X(2), Y(2), Z(2),
	A1(2), B1(2), C1(2), D1(2), E1(2), F1(2), G1(2), S, Rout(2));
	Mux_32_a_18Bits_3: Mux32_a_1 port map (A(3), B(3), C(3), D(3), E(3), F(3), G(3), H(3), I(3), J(3),
	K(3), L(3), M(3), N(3), O(3), P(3), Q(3), R(3), Si(3), T(3), U(3), W(3), X(3), Y(3), Z(3),
	A1(3), B1(3), C1(3), D1(3), E1(3), F1(3), G1(3), S, Rout(3));
	Mux_32_a_18Bits_4: Mux32_a_1 port map (A(4), B(4), C(4), D(4), E(4), F(4), G(4), H(4), I(4), J(4),
	K(4), L(4), M(4), N(4), O(4), P(4), Q(4), R(4), Si(4), T(4), U(4), W(4), X(4), Y(4), Z(4),
	A1(4), B1(4), C1(4), D1(4), E1(4), F1(4), G1(4), S, Rout(4));
	Mux_32_a_18Bits_5: Mux32_a_1 port map (A(5), B(5), C(5), D(5), E(5), F(5), G(5), H(5), I(5), J(5),
	K(5), L(5), M(5), N(5), O(5), P(5), Q(5), R(5), Si(5), T(5), U(5), W(5), X(5), Y(5), Z(5),
	A1(5), B1(5), C1(5), D1(5), E1(5), F1(5), G1(5), S, Rout(5));
	Mux_32_a_18Bits_6: Mux32_a_1 port map (A(6), B(6), C(6), D(6), E(6), F(6), G(6), H(6), I(6), J(6),
	K(6), L(6), M(6), N(6), O(6), P(6), Q(6), R(6), Si(6), T(6), U(6), W(6), X(6), Y(6), Z(6),
	A1(6), B1(6), C1(6), D1(6), E1(6), F1(6), G1(6), S, Rout(6));
	Mux_32_a_18Bits_7: Mux32_a_1 port map (A(7), B(7), C(7), D(7), E(7), F(7), G(7), H(7), I(7), J(7),
	K(7), L(7), M(7), N(7), O(7), P(7), Q(7), R(7), Si(7), T(7), U(7), W(7), X(7), Y(7), Z(7),
	A1(7), B1(7), C1(7), D1(7), E1(7), F1(7), G1(7), S, Rout(7));
	
	Mux_32_a_18Bits_8: Mux32_a_1 port map (A(8), B(8), C(8), D(8), E(8), F(8), G(8), H(8), I(8), J(8),
	K(8), L(8), M(8), N(8), O(8), P(8), Q(8), R(8), Si(8), T(8), U(8), W(8), X(8), Y(8), Z(8),
	A1(8), B1(8), C1(8), D1(8), E1(8), F1(8), G1(8), S, Rout(8));
	Mux_32_a_18Bits_9: Mux32_a_1 port map (A(9), B(9), C(9), D(9), E(9), F(9), G(9), H(9), I(9), J(9),
	K(9), L(9), M(9), N(9), O(9), P(9), Q(9), R(9), Si(9), T(9), U(9), W(9), X(9), Y(9), Z(9),
	A1(9), B1(9), C1(9), D1(9), E1(9), F1(9), G1(9), S, Rout(9));
	Mux_32_a_18Bits_10: Mux32_a_1 port map (A(10), B(10), C(10), D(10), E(10), F(10), G(10), H(10), I(10), J(10),
	K(10), L(10), M(10), N(10), O(10), P(10), Q(10), R(10), Si(10), T(10), U(10), W(10), X(10), Y(10), Z(10),
	A1(10), B1(10), C1(10), D1(10), E1(10), F1(10), G1(10), S, Rout(10));
	Mux_32_a_18Bits_11: Mux32_a_1 port map (A(11), B(11), C(11), D(11), E(11), F(11), G(11), H(11), I(11), J(11),
	K(11), L(11), M(11), N(11), O(11), P(11), Q(11), R(11), Si(11), T(11), U(11), W(11), X(11), Y(11), Z(11),
	A1(11), B1(11), C1(11), D1(11), E1(11), F1(11), G1(11), S, Rout(11));
	Mux_32_a_18Bits_12: Mux32_a_1 port map (A(12), B(12), C(12), D(12), E(12), F(12), G(12), H(12), I(12), J(12),
	K(12), L(12), M(12), N(12), O(12), P(12), Q(12), R(12), Si(12), T(12), U(12), W(12), X(12), Y(12), Z(12),
	A1(12), B1(12), C1(12), D1(12), E1(12), F1(12), G1(12), S, Rout(12));
	Mux_32_a_18Bits_13: Mux32_a_1 port map (A(13), B(13), C(13), D(13), E(13), F(13), G(13), H(13), I(13), J(13),
	K(13), L(13), M(13), N(13), O(13), P(13), Q(13), R(13), Si(13), T(13), U(13), W(13), X(13), Y(13), Z(13),
	A1(13), B1(13), C1(13), D1(13), E1(13), F1(13), G1(13), S, Rout(13));
	Mux_32_a_18Bits_14: Mux32_a_1 port map (A(14), B(14), C(14), D(14), E(14), F(14), G(14), H(14), I(14), J(14),
	K(14), L(14), M(14), N(14), O(14), P(14), Q(14), R(14), Si(14), T(14), U(14), W(14), X(14), Y(14), Z(14),
	A1(14), B1(14), C1(14), D1(14), E1(14), F1(14), G1(14), S, Rout(14));
	Mux_32_a_18Bits_15: Mux32_a_1 port map (A(15), B(15), C(15), D(15), E(15), F(15), G(15), H(15), I(15), J(15),
	K(15), L(15), M(15), N(15), O(15), P(15), Q(15), R(15), Si(15), T(15), U(15), W(15), X(15), Y(15), Z(15),
	A1(15), B1(15), C1(15), D1(15), E1(15), F1(15), G1(15), S, Rout(15));
	
	Mux_32_a_18Bits_16: Mux32_a_1 port map (A(16), B(16), C(16), D(16), E(16), F(16), G(16), H(16), I(16), J(16),
	K(16), L(16), M(16), N(16), O(16), P(16), Q(16), R(16), Si(16), T(16), U(16), W(16), X(16), Y(16), Z(16),
	A1(16), B1(16), C1(16), D1(16), E1(16), F1(16), G1(16), S, Rout(16));
	Mux_32_a_18Bits_17: Mux32_a_1 port map (A(17), B(17), C(17), D(17), E(17), F(17), G(17), H(17), I(17), J(17),
	K(17), L(17), M(17), N(17), O(17), P(17), Q(17), R(17), Si(17), T(17), U(17), W(17), X(17), Y(17), Z(17),
	A1(17), B1(17), C1(17), D1(17), E1(17), F1(17), G1(17), S, Rout(17));
	Mux_32_a_18Bits_18: Mux32_a_1 port map (A(18), B(18), C(18), D(18), E(18), F(18), G(18), H(18), I(18), J(18),
	K(18), L(18), M(18), N(18), O(18), P(18), Q(18), R(18), Si(18), T(18), U(18), W(18), X(18), Y(18), Z(18),
	A1(18), B1(18), C1(18), D1(18), E1(18), F1(18), G1(18), S, Rout(18));
	Mux_32_a_18Bits_19: Mux32_a_1 port map (A(19), B(19), C(19), D(19), E(19), F(19), G(19), H(19), I(19), J(19),
	K(19), L(19), M(19), N(19), O(19), P(19), Q(19), R(19), Si(19), T(19), U(19), W(19), X(19), Y(19), Z(19),
	A1(19), B1(19), C1(19), D1(19), E1(19), F1(19), G1(19), S, Rout(19));
	Mux_32_a_18Bits_20: Mux32_a_1 port map (A(20), B(20), C(20), D(20), E(20), F(20), G(20), H(20), I(20), J(20),
	K(20), L(20), M(20), N(20), O(20), P(20), Q(20), R(20), Si(20), T(20), U(20), W(20), X(20), Y(20), Z(20),
	A1(20), B1(20), C1(20), D1(20), E1(20), F1(20), G1(20), S, Rout(20));

end Mux_32_a_1_21Bits;