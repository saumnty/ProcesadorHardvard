library IEEE;
use IEEE.std_logic_1164.all;

entity Procesador_Test is
end Procesador_Test;

architecture Procesador_Test of Procesador_Test is

component Procesador is
	port(
	clk: in std_logic;
	Mem_Codigos_Data: out std_logic_vector (20 downto 0);
	DCout, DAout, DBout: out std_logic_vector (2 downto 0);
	WIRout, WCWout: out std_logic;
	Wout, WEout, Miout, MMout, MWout: out std_logic;	
	MBout, MCout, WPCout: out std_logic;
	Selc_out: out std_logic_vector(4 downto 0);
	Carry_out,Vo_out,Zero_out,Signo_out: out std_logic;
	J_Result, Sv_result: out std_logic;
	PCout: out std_logic_vector (7 downto 0);
	Result: out std_logic_vector (7 downto 0));
end component;

signal clk: std_logic;
signal MWC: std_logic := '1';
signal Mem_Codigos_Data: std_logic_vector (20 downto 0);
signal DCout, DAout, DBout: std_logic_vector (2 downto 0);
signal WIRout, WCWout: std_logic;
signal Wout, WEout, Miout, MMout, MWout: std_logic;
signal MBout, MCout, WPCout: std_logic;
signal Selc_out: std_logic_vector (4 downto 0);
signal Carry_out,Vo_out,Zero_out,Signo_out: std_logic;
signal J_Result, Sv_result: std_logic;
signal PCout: std_logic_vector (7 downto 0);
signal Result: std_logic_vector (7 downto 0);

begin

Procesador_F: Procesador port map(clk, Mem_Codigos_Data, DCout, DAout, DBout, WIRout, WCWout, Wout, WEout,
Miout, MMout, MWout, MBout, MCout, WPCout, Selc_out, Carry_out, Vo_out, Zero_out, Signo_out, J_Result, Sv_result, PCout, Result);

process is
	begin
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait for 4 ns;
	clk <= '0';
	wait for 4 ns;
	clk <= '1';
	wait;
end process;
end Procesador_Test;